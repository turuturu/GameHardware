
/*
Video sync generator, used to drive a simulated CRT.
To use:
- Wire the hsync and vsync signals to top level outputs
- Add a 3-bit (or more) "rgb" output to the top level
*/

module hvsync_generator #(
  parameter H_DISPLAY       = 256, // horizontal display width // 640
  parameter H_BACK          =  23, // horizontal left border (back porch) // 48
  parameter H_FRONT         =   7, // horizontal right border (front porch) // 16
  parameter H_SYNC          =  23, // horizontal sync width // 96
  // vertical constants
  parameter V_DISPLAY       = 240, // vertical display height // 480
  parameter V_TOP           =   5, // vertical top border // 33
  parameter V_BOTTOM        =  14, // vertical bottom border // 10
  parameter V_SYNC          =   3, // vertical sync # lines // 2
  parameter DATA_WIDTH      =   10
)
(
  input clk,
  input reset,
  output reg hsync, vsync,
  output display_on,
  output reg [DATA_WIDTH-1:0] hpos,
  output reg [DATA_WIDTH-1:0] vpos
);

  // declarations for TV-simulator sync parameters
  // horizontal constants
  // derived constants
  parameter H_SYNC_START    = H_DISPLAY + H_FRONT;
  parameter H_SYNC_END      = H_DISPLAY + H_FRONT + H_SYNC - 1;
  parameter H_MAX           = H_DISPLAY + H_BACK + H_FRONT + H_SYNC - 1;
  parameter V_SYNC_START    = V_DISPLAY + V_BOTTOM;
  parameter V_SYNC_END      = V_DISPLAY + V_BOTTOM + V_SYNC - 1;
  parameter V_MAX           = V_DISPLAY + V_TOP + V_BOTTOM + V_SYNC - 1;

  wire hmaxxed = (hpos == H_MAX) || reset;	// set when hpos is maximum
  wire vmaxxed = (vpos == V_MAX) || reset;	// set when vpos is maximum
  
  // horizontal position counter
  always @(posedge clk)
  begin
    hsync <= ~(hpos>=H_SYNC_START && hpos<=H_SYNC_END);
    if(hmaxxed)
      hpos <= 0;
    else
      hpos <= hpos + 1;
  end

  // vertical position counter
  always @(posedge clk)
  begin
    vsync <= ~(vpos>=V_SYNC_START && vpos<=V_SYNC_END);
    if(hmaxxed)
      if (vmaxxed)
        vpos <= 0;
      else
        vpos <= vpos + 1;
  end
  
  // display_on is set when beam is in "safe" visible frame
  assign display_on = (hpos<H_DISPLAY) && (vpos<V_DISPLAY);

endmodule
